* NGSPICE file created from posoco2000.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

.subckt posoco2000 clk segm[0] segm[1] segm[2] segm[3] segm[4] segm[5] segm[6] segm[7]
+ sel[0] sel[1] sel[2] sel[3] sel[4] sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__163__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_131_ net16 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_114_ net8 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__126__A2 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__077__I _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput7 net7 sel[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_130_ _072_ _048_ _070_ _042_ _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__153__CLK clknet_1_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output12_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_113_ _058_ _051_ _060_ _044_ _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput8 net8 sel[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput10 net10 sel[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__088__I dut.count\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output2_I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__135__B _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__096__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__147__A1 _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__138__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_112_ _059_ _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__166__CLK clknet_1_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput9 net9 sel[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput11 net11 sel[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__099__I _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__135__C net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__138__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_111_ _038_ _031_ _054_ _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput12 net12 sel[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__156__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__101__B1 _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_110_ net9 _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output10_I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput13 net13 sel[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__101__B2 _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__169__CLK clknet_1_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_169_ _017_ clknet_1_0__leaf_clk dut.count\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xposoco2000_17 segm[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput14 net14 sel[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__102__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__154__D _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__101__A2 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__110__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__105__I dut.count\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_168_ _016_ clknet_1_1__leaf_clk dut.count\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__162__D _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_099_ _047_ _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xposoco2000_18 segm[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__157__D _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__159__CLK clknet_1_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput15 net15 sel[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__094__B dut.count\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__108__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__165__D _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_167_ _015_ clknet_1_1__leaf_clk dut.count\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_098_ net12 _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__116__I _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__140__A1 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput16 net16 sel[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__122__A1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_clk clk clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__168__D _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__113__B2 _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__119__I dut.count\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_166_ _014_ clknet_1_0__leaf_clk net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_097_ _042_ _044_ _046_ _048_ _049_ _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_149_ _028_ _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__113__A2 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output9_I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_165_ _013_ clknet_1_0__leaf_clk net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_096_ net13 _049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_148_ _021_ _074_ _027_ _028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_079_ dut.count\[1\] _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__151__I _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_164_ _012_ clknet_1_0__leaf_clk net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__146__I _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_095_ _047_ _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__143__A1 _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_078_ _031_ _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_147_ _032_ _039_ _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__149__I _028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__162__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_163_ _011_ clknet_1_1__leaf_clk net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_094_ dut.count\[1\] dut.count\[2\] dut.count\[3\] _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_146_ _026_ _017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_077_ _030_ _031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_129_ net15 _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output7_I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__152__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_162_ _010_ clknet_1_1__leaf_clk net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_093_ _045_ _035_ _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_clk_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_145_ _035_ _025_ _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_076_ dut.count\[3\] _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__122__B net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__083__I _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_128_ _066_ _071_ _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_161_ _009_ clknet_1_1__leaf_clk net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_092_ _030_ _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__128__A1 _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_144_ _032_ _069_ _065_ _025_ _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__165__CLK clknet_1_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__133__B _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_127_ net3 _062_ _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__082__A1 _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_160_ _008_ clknet_1_0__leaf_clk net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__137__A2 _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_091_ _043_ _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_143_ _015_ _043_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_126_ _046_ _065_ _066_ _068_ _070_ _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__144__B _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_109_ _015_ _044_ _056_ _048_ _057_ _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__155__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output5_I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_090_ _033_ _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_142_ _065_ _023_ _024_ _040_ _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_23_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_125_ _037_ _069_ _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_108_ net10 _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__168__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_141_ net5 _047_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_124_ _033_ _054_ _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_107_ _055_ _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__100__A2 _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__094__A1 dut.count\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__085__A1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__152__D _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_140_ _040_ _022_ _023_ _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__158__CLK clknet_1_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output13_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_123_ _055_ _067_ _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__103__B1 _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__160__D _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_106_ _030_ _054_ _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__155__D _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__094__A2 dut.count\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__085__A2 dut.count\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output3_I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__087__B _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__163__D _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__130__B2 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_122_ _038_ _064_ _031_ net6 _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__158__D _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__103__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_105_ dut.count\[2\] _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__097__B1 _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__114__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__171__D _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__085__A3 dut.count\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__166__D _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__130__A2 _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__117__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_121_ _064_ _059_ _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_1_0__f_clk clknet_0_clk clknet_1_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__103__A2 _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_104_ dut.count\[0\] _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__097__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__115__B1 _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_120_ _038_ _064_ _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__103__A3 _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__171__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output11_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_103_ _042_ _034_ _046_ _048_ _053_ _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__097__A2 _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__142__A1 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__142__B2 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output1_I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__115__B2 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__106__A1 _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_102_ net11 _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__097__A3 _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__139__I _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__161__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__133__A2 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__115__A2 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_101_ _050_ _051_ _052_ _046_ _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_24_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__118__B1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__109__B1 _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_100_ _041_ _044_ _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__081__I dut.count\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__076__I dut.count\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__127__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__118__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__118__B2 _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__109__A1 _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__164__CLK clknet_1_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__084__I dut.count\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_159_ _007_ clknet_1_0__leaf_clk net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__079__I dut.count\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__092__I _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__127__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__118__A2 _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__109__A2 _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_158_ _006_ clknet_1_0__leaf_clk net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_089_ _041_ _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__095__I _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__154__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_1__f_clk clknet_0_clk clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__118__A3 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__109__A3 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__098__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_157_ _005_ clknet_1_0__leaf_clk net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_088_ dut.count\[0\] _041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__167__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_156_ _004_ clknet_1_1__leaf_clk net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_087_ _032_ _036_ _040_ _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_139_ _075_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__148__A2 _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output8_I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__157__CLK clknet_1_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_155_ _003_ clknet_1_1__leaf_clk net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_086_ _037_ _039_ _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_138_ net2 _062_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__082__B net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__153__D _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_171_ _019_ clknet_1_1__leaf_clk net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__120__A1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__111__A1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_154_ _002_ clknet_1_1__leaf_clk net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_085_ _038_ dut.count\[1\] dut.count\[2\] _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_18_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__104__I dut.count\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_137_ _060_ _075_ _020_ _021_ _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__161__D _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__156__D _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput1 net1 segm[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_170_ _018_ clknet_1_1__leaf_clk dut.count\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__164__D _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_153_ _001_ clknet_1_0__leaf_clk net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_084_ dut.count\[0\] _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__159__D _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__087__A1 _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_136_ _037_ _039_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_119_ dut.count\[1\] _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__150__B1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__167__D _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput2 net2 segm[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output6_I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_152_ _000_ clknet_1_1__leaf_clk net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_083_ _030_ _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__170__CLK clknet_1_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_135_ _064_ _035_ _032_ net1 _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__131__I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_118_ _042_ _034_ _056_ _062_ _063_ _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__150__B2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__141__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput3 net3 segm[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_151_ _029_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_082_ _034_ _035_ net14 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__129__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_134_ _033_ _054_ _031_ _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__160__CLK clknet_1_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_117_ net7 _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__150__A2 _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__141__A2 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput4 net4 segm[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_150_ _041_ _034_ _056_ _062_ net4 _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_27_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_081_ dut.count\[2\] _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_133_ _073_ _051_ _074_ _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_116_ _047_ _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__150__A3 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__126__B1 _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput5 net5 segm[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output4_I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_080_ _033_ _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_132_ _041_ _037_ _069_ _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_115_ _061_ _051_ _052_ _056_ _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__144__A1 _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__126__A1 _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput6 net6 segm[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

