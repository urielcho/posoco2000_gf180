magic
tech gf180mcuC
magscale 1 5
timestamp 1670198804
<< obsm1 >>
rect 672 1538 29288 28254
<< metal2 >>
rect 1344 29600 1400 29900
rect 7728 29600 7784 29900
rect 14112 29600 14168 29900
rect 20496 29600 20552 29900
rect 26880 29600 26936 29900
rect 0 100 56 400
rect 6048 100 6104 400
rect 12432 100 12488 400
rect 18816 100 18872 400
rect 25200 100 25256 400
<< obsm2 >>
rect 14 29570 1314 29600
rect 1430 29570 7698 29600
rect 7814 29570 14082 29600
rect 14198 29570 20466 29600
rect 20582 29570 26850 29600
rect 26966 29570 29106 29600
rect 14 430 29106 29570
rect 86 400 6018 430
rect 6134 400 12402 430
rect 12518 400 18786 430
rect 18902 400 25170 430
rect 25286 400 29106 430
<< metal3 >>
rect 29600 26880 29900 26936
rect 100 25200 400 25256
rect 29600 20496 29900 20552
rect 100 18816 400 18872
rect 29600 14112 29900 14168
rect 100 12432 400 12488
rect 29600 7728 29900 7784
rect 100 6048 400 6104
rect 29600 1344 29900 1400
<< obsm3 >>
rect 9 26966 29600 28238
rect 9 26850 29570 26966
rect 9 25286 29600 26850
rect 9 25170 70 25286
rect 430 25170 29600 25286
rect 9 20582 29600 25170
rect 9 20466 29570 20582
rect 9 18902 29600 20466
rect 9 18786 70 18902
rect 430 18786 29600 18902
rect 9 14198 29600 18786
rect 9 14082 29570 14198
rect 9 12518 29600 14082
rect 9 12402 70 12518
rect 430 12402 29600 12518
rect 9 7814 29600 12402
rect 9 7698 29570 7814
rect 9 6134 29600 7698
rect 9 6018 70 6134
rect 430 6018 29600 6134
rect 9 1430 29600 6018
rect 9 1314 29570 1430
rect 9 910 29600 1314
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
rect 25264 1538 25424 28254
<< obsm4 >>
rect 19222 7009 19250 7439
<< labels >>
rlabel metal3 s 29600 1344 29900 1400 6 clk
port 1 nsew signal input
rlabel metal3 s 29600 7728 29900 7784 6 segm[0]
port 2 nsew signal output
rlabel metal2 s 18816 100 18872 400 6 segm[1]
port 3 nsew signal output
rlabel metal3 s 29600 20496 29900 20552 6 segm[2]
port 4 nsew signal output
rlabel metal3 s 29600 26880 29900 26936 6 segm[3]
port 5 nsew signal output
rlabel metal3 s 100 25200 400 25256 6 segm[4]
port 6 nsew signal output
rlabel metal2 s 20496 29600 20552 29900 6 segm[5]
port 7 nsew signal output
rlabel metal2 s 0 100 56 400 6 segm[6]
port 8 nsew signal output
rlabel metal2 s 7728 29600 7784 29900 6 segm[7]
port 9 nsew signal output
rlabel metal2 s 25200 100 25256 400 6 sel[0]
port 10 nsew signal output
rlabel metal2 s 6048 100 6104 400 6 sel[1]
port 11 nsew signal output
rlabel metal2 s 14112 29600 14168 29900 6 sel[2]
port 12 nsew signal output
rlabel metal3 s 100 6048 400 6104 6 sel[3]
port 13 nsew signal output
rlabel metal3 s 100 12432 400 12488 6 sel[4]
port 14 nsew signal output
rlabel metal2 s 26880 29600 26936 29900 6 sel[5]
port 15 nsew signal output
rlabel metal2 s 12432 100 12488 400 6 sel[6]
port 16 nsew signal output
rlabel metal3 s 100 18816 400 18872 6 sel[7]
port 17 nsew signal output
rlabel metal2 s 1344 29600 1400 29900 6 sel[8]
port 18 nsew signal output
rlabel metal3 s 29600 14112 29900 14168 6 sel[9]
port 19 nsew signal output
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 20 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 20 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 21 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 28254 6 vss
port 21 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 663342
string GDS_FILE /home/urielcho/Proyectos_caravel/gf180nm/posoco2000/openlane/posoco2000/runs/22_12_04_18_05/results/signoff/posoco2000.magic.gds
string GDS_START 135582
<< end >>

